1 10 11 100 101 110 111 1000 1001 1010 1011 1100 1101 1110 1111 10000 10001 10010 10011 10100 10101 10110 10111 11000 11001 11010 11011 11100 11101 11110 11111 100000 11111 11110 1101 11001 11000 10111 10110 10101 10100 10011 10010 10001 10000 1111 1110 1101 1100 1011 1010 1001 1000 111 110 101 100 11 10 1 0 10001001 10001100 10001101 10001111 10010000 10010001 10010010 10010011 10010100 10010101 10010110 10010111 10011000 10011001 10011010 10011011 10011100 10011101 10011110 10011111 10100001 10100010 10100011 10100100 10100101 10100110 10100111 10101000 10101001 10101010 10101011 10101100 10101101 10101110 10101111 10110000 10111000 10111001 10111010 10111011 10111100 10111101 10111110 10111111 11000000 11000001 11000010 11000011 11000100 11000101 11000110 11000111 11001000 11001001 11001010 11001011 11001100 11001101 11001110 11001111 11010000 11010001 11010010 11010011 11010100 11010101 11010110 11010111 11011000 11011001 11011010 11011011 11011100 11011101 11011110 11011111 11100000 11100001 11100010 11100011 11100100 11100101 11100110 11100111 11101000 11101001 11101010 11101011 11101100 11101101 11101110 11101111 11110000 11110001 11110010 11110011 11110100 11110101 11110110 11110111 11111000 11111001 11111010 11111011 11111100 11111101 11111110 11111111 11111110 11110111 11110110 11110101 11110100 11110011 11110010 11110001 11110000 11101110 11101101 11101100 11101011 11101010 11101001 11101000 11100111 11100110 11100101 11100100 11100011 11100001 11100000 11011110 11011101 11011100 11011011 11011010 11011001 11011000 11010111 11010110 11010101 11010100 11010011 11010010 11010001 11010000 11001111 11001110 11000111 11000110 11000101 11000100 11000011 11000010 11000001 11000000 10111110 10011111 10011110 10001111 10001110 10001111 10000110 10000101 10000100 10000011 10000010 10000001 10000000 01111111 01111110 00111111 00111110 00011111 00011110 00001111 00001110 00001101 00001100 00001011 00001010 00001001 00001000 00000110 00000010 0 1 2 10 11 12 20 21 22 100 101 102 110 111 112 120 121 122 200 201 202 210 211 212 220 221 222 1000 1001 1002 1010 1011 1012 1020 1021 1022 1100 1101 1102 1110 1111 1112 1120 1121 1122 1200 1201 1202 1210 1211 1212 1220 1221 1222 2000 2001 2002 2010 2011 2012 2020 2021 2022 2100 2101 2102 2110 2111 2112 2120 2121 2122 2200 2201 2202 2210 2211 2212 2220 2221 2222 10000 10001 10002 10010 10011 10021 10022 10100 10101 10102 10110 10111 10112 10120 10121 10122 10200 10201 10220 10210 10211 10212 10220 10221 10222 11000 11100 11101 11102 11110 11111 11112 11120 11121 11122 11200 11202 11210 11211 11212 11220 11221 11222 12000 12001 12002 12010 12011 12012 12020 12021 12022 12100 12101 12102 12110 12111 12112 12120 12121 12122 12200 12202 12210 12211 12212 12220 12221 12222 20000 20001 20002 200010 20001 20002 20010 20011 20012 20020 20021 20022 20100 20101 20102 20110 20111 20112 20120 20121 20122 20200 20201 20202 20210 20211 20212 20220 20221 20222 21000 21001 21002 21012 21020 21021 21022 21100 21101 21102 21110 21111 21112 21120 21121 21122 21200 21201 21202 21210 21211 21212 21220 21221 21222 22000 22001 22002 22002 22010 22012 22020 22021 22022 22100 22102 22110 22111 22112 22120 22121 22122 22200 22201 22202 22210 22211 22212 22220 22221 22222 100000 100001 100002 100010 100011 100012 100020 100021 100022 100100 100102 100110 100111 100112 100120 100121 100122 100200 100202 100210 100211 100212 100220 100221 100222 101000 101001 101002 101010 101011 101012 101020 101021 101022 101100 101102 101110 101111 101112 101120 101121 101122 101200 101201 101202 101210 101211 101212 101220 101221 101222 102000 102001 102002 102010 102011 102012 102020 102021 102022 102100 102101 102102 102110 102111 102112 102120 102121 102122 102200 102201 102202 102210 102211 102212 102220 102221 102222 110000 110001 110002 110010 110011 110012 110020 110021 110022 110100 110101 110102 110110 110111 110112 110120 110121 110122 110200 110201 110202 110210 110211 110212 110220 110221 110222 111000 111001 111002 111010 111011 111012 111020 111021 111022 111100 111101 111102 111110 111111 111112 111120 111121 111122 111200 111201 111202 111210 111211 111212 111220 111221 111222 112000 112001 112002 112010 112011 112012 112020 112021 112022 112100 112101 112102 112110 112111 112112 112120 112121 112122 112200 112201 112202 112210 112212 112220 112221 112222 120000 120001 120002 120010 120011 120012 100222 120021 120022 120100 120101 120102 120110 120111 120112 120120 120121 120122 120200 120201 120202 120210 120211 120212 120220 120221 120222 121000 121001 121002 121010 121011 121012 121020 121201 121022 121100 121101 121102 121110 121111 121112 121120 121121 121122 121200 121201 121202 121210 121211 121212 121220 121221 121222 122000 122001 122002 122010 122011 122012 122020 122021 122022 122100 122101 122102 122110 122111 122112 122120 122121 122122 122200 122201 122202 122210 122211 122212 122220 122221 122222 200000 200001 200002 200010 200011 200012 200020 200021 200022 200100 200101 200102 200110 200111 200112 200120 200121 200122 200200 200202 200210 200211 200212 200220 200221 200222 201000 201001 201002 201010 201011 201012 201020 201021 201022 201100 201101 201102 201110 201111 201112 201120 201121 201122 201200 201201 201202 201210 201211 201212 201220 201221 201222 202000 202001 202002 202010 202011 202012 202020 202021 202022 202100 202101 202102 202110 202111 202112 202120 202121 202122 202200 202202 202210 202211 202212 202220 202221 202222 210000 210001 210002 210010 210011 210012 210020 210021 210022 210100 210101 210102 210110 210111 210112 210120 210121 210122 210200 210201 210202 210210 210211 210212 210220 210221 210222 211000 211001 211002 211010 211011 211012 211020 211021 211022 211100 211101 211102 211110 211111 211112 211120 211121 211122 211200 211201 211202 211210 211211 211212 211220 211221 211222 212000 212001 212002 212011 212012 212020 212021 210221 212022 212100 212101 212102 212110 212111 212112 212120 212121 212122 212200 212201 212202 212210 212211 212212 212220 212221 212222 220000 220001 220002 220010 220011 220012 220020 220021 220022 220100 220101 220102 220110 220111 220112 220120 220121 220122 220200 220201 220202 220210 220211 220212 220220 220221 220222 221000 221001 221002 221010 221011 221012 221020 221021 221022 221100 221101 221102 221110 221111 221112 221120 221121 221122 221200 221201 221202 221210 221211 221212 221220 221221 221222 222000 222001 222002 222010 222011 222012 222020 222021 222022 222100 222101 222102 222110 222111 222112 222120 222121 222122 222200 222201 222202 222210 222211 222212 222220 222221 222222 1000000 1000001 1000002 1000010 100011 100012 1000011 1000012 1000020 1000021 1000022 1000100 1000101 1000102 1000110 1000111 1000112 1000120 1000121 1000122 1000200 1000201 1000202 1000210 1000211 1000212 1000220 1000221 1000222 1001000 1001001 1001002 1001010 1001011 1001012 1001020 1001021 1002000 1002001 1002002 1002001 1002010 1002012 1002020 1002021 1002022 1002100 1002101 1002102 1002110 1002111 1002112 1002120 1002121 1002122 1002200 1002201 1002202 1002210 1002211 1002212 1002220 1002221 1002222 1010000 1010001 1010002 1010010 1010011 1010012 1010020 1010021 1010022 1010100 1010101 1010102 1010110 1010111 1010112 1010120 1010121 1010122 1010200 1010201 1010202 1010210 1010212 1010220 1010221 1010222 1011000 1011001 1011002 1011010 1011011 1011012 1011020 1011021 1011022 1011100 1011102 1011110 1011111 1011112 1011120 1011121 1011122 1011200 1011201 1011202 1011210 1011211 1011212 1011220 1011221 1011222 1012000 1012001 1012002 1012010 1012011 1012012 1012020 1012021 1012022 1012100 1012101 1012102 1201 1012112 1012120 1012121 1012122 101200 1012200 1012201 1012202 1012210 1012211 1012212 1012220 1012221 1012222 1020000 1020001 1020002 1020010 1020011 1020012 1020020 1020021 1020022 1020100 1020101 1020101 1020102 1020110 1020112 1020120 1020121 1020122 1020200 1020201 1020202 1020210 1020211 1020212 1020220 1020221 1020222 1021000 1021001 1021002 1021010 1021011 1021012 1021020 1021021 1021022 1021100 1021110 1021102 1021111 1021112 1021120 1021121 1021122 1021200 1021201 1021202 1021210 1021211 1021212 1021220 1201212 1021220 1021221 1021222 1022000 1022001 1022002 1022010 1022011 1022012 1022020 1022021 1022022 1022100 1022101 1022102 1022110 1022111 1022112 1022120 1022121 1022122 1022200 1022201 1022202 1022210 1022211 1022212 1022220 1022221 1022222 1100000 1100002 1100010 1100011 1100012 1100020 1100021 1100022 1100100 1100101 1100102 1100110 1100111 1100112 1100120 1100121 1100122 1100200 1100201 1100202 1100210 1100211 1100212 1100220 1100221 1100222 1101000 1101001 1101002 1101010 1101011 1101012 1101020 1101021 1101022 1101100 1101101 1101102 1101110 1101111 1101112 1101120 1101122 1101200 1101201 1101202 1101210 1101211 1101212 1101220 1101221 1101222 1102000 1102001 1102002 1102010 1102011 1102012 1102020 1102021 1102022 1102100 1102101 1102102 1102111 1102112 1102120 1102121 1102122 1102200 1102220 1102221 1102222 1110000 1110001 1110002 1110010 1110011 1110012 1110020 1110021 1110022 1110100 1111010 1110101 1110102 1110110 1110111 1110112 1110120 1110121 1110122 1110200 1110201 1110202 1110210 1110211 1110212 1110220 1110221 1110222 1111000 1111001 1111002 1111010 1111100 1111001 1111110 1111111 1111112 1111120 1111200 1111201 1111202 1111210 1112000 1112001 1112002 1112010 1112011 1112012 1112020 1112021 1112022 1112100 1112101 1112102 1112110 1112111 1112112 1112120 1112121 1112122 1112200 1112201 1112202 1112210 1112211 1112212 1112220 1112221 1112222 1120000 1120001 1120002 1120010 1120011 1120012 1120020 1120021 1120022 1120100 1120101 1120200 1120201 1120202 1120210 1120211 1120212 1120220 1120221 1120222 1121000 1121001 1121002 1121010 1121011 1121012 1121020 1121021 1121022 1121100 1121110 1121111 1121112 1121120 1121121 1121122 1121200 1121201 1121202 1121210 1121211 1121212 1121220 1121221 1121222 1122000 1122001 1122002 1122010 1122011 1122012 1122020 1122021 1122022 1122100 1122101 1122102 1122110 1122111 1122112 1122120 1122121 1122122 1122200 1122201 1122202 1122210 1122211 1122212 1122220 1122221 1122222 1200000 1200001 1200002 1200010 1200011 1200012 1200020 1200021 1200022 1200100 1200101 1200102 1200110 1200111 1200112 1200120 1200121 1200122 1200200 1200201 1200202 1200210 1200211 1200212 1200220 1200221 1200222 1201000 1201001 1201002 1201010 1201011 1201012 1201012 1201021 1201022 1201100 1201101 1201102 1201110 1201111 1201112 1201120 1201121 1201122 1201200 1201201 1201202 1201210 1201211 1201212 1201220 1201222 1202000 1202001 1202002 1202010 1202011 1202012 1202020 1202021 1202022 1202100 1202101 1202102 1202110 1202111 1202112 1202120 1202121 1202122 1202200 1202201 1202202 1202210 1202211 1202212 1202220 1202221 1202222 1210000 1210001 1210002 1210010 1210011 1210012 1210020 1210021 1210022 1210100 1201101 1210121 1210122 1211000 1211001 1211002 1211010 1211011 1211012 1211020 1211021 1211022 1211100 1211101 1211102 1211110 1211111 1211112 1211120 1211121 1211112 1211200 1211201 1211202 1211210 1211212 1211220 1211212 1211220 1211221 1211222 1212000 1212001 1212002 1212010 1212011 1212012 1212020 1212021 1212022 1212100 1212101 1212102 1212110 1212111 1212112 1212120 1212121 1212122 1212200 1212201 1212202 1212210 1212211 1212212 1212220 1212221 1212222 1220000 1220001 1220002 1220010 1220011 1220012 1220020 1220021 1220022 1220100 1220101 1220102 1220110 1220111 1220112 1220120 1220121 1220122 1220200 1220201 1220202 1220210 1220211 1220212 1220220 1220221 1220222 1221000 1221001 1221002 1221010 1221011 1221012 1221020 1221021 1221022 1221100 1221101 1221102 1221110 1221111 1221112 1221120 1221121 1221122 1221200 1221201 1221202 1221210 1221211 1221212 1221220 1221221 1221222 1222000 1222001 1222002 1222010 1222011 1222012 1222020 1222021 1222022 1222100 1222101 1222102 1222110 1222111 1222112 1222120 1222121 1222122 1222200 1222201 1222202 1222210 1222211 1222212 1222220 1222221 1222222 2000000 2000001 2000002 2000010 2000011 2000012 2000020 2000021 2000002 2000022 2000100 2000101 2000102 2000110 2000111 2000112 2000120 2000121 2000122 2000200 2000201 2000202 2000210 2000211 2000212 2000220 2000221 2000222 2001000 2001001 2001002 2001010 2001011 2001012 2001020 2001021 2001022 2001100 2001101 2001102 2001110 2001111 2001112 2001120 2001121 2001122 2001200 2001201 2001202 2001210 2001211 2001212 2001220 2001221 2001222 2002000 2002001 2002002 2002010 2002011 2002012 2002020 2002021 2002022 2002100 2002101 2002102 2002110 2002111 2002112 2002120 2002121 2002122 2002200 2002201 2002202 2002210 2002211 2002212 2002220 2002221 2002222 2010000 2010002 2010010 2010011 2010012 2010020 2010021 2010022 2010100 2010101 2010102 2010110 2010111 2010120 2010121 2010122 2010200 2010201 2010202 2010201 2010200 2010122 2010121 2010120 2010110 2010102 2010101 2010100 2010022 2010021 2010020 2010012 2010011 2010010 2010002 2010001 2010000 2002222 2002202 2002201 2002200 2002122 2002121 2002120 2002112 2002111 2002110 2002102 2002101 2002100 2002022 2002021 2002020 2002012 2002011 2002010 2000200 2000122 2000121 2000120 2000112 2000111 2000110 2000102 2000101 2000100 2000022 2000021 2000020 2000012 2000011 2000010 2000002 2000001 2000000 1222222 1212222 1220000 1210222 1210221 1210220 1210212 1210211 1210210 1210202 1210201 1210200 1210122 1210121 1210120 1210112 1210111 1210110 1210102 1210101 1210100 1210022 1210021 1210020 1210012 1210011 1210010 1210002 1210001 1210000 1202222 1202221 1202220 1202212 1202211 1202210 1202202 1202201 1202200 1202122 1202121 1202120 1202112 1202111 1202110 1202102 1202101 1202100 1202100 1202022 1202021 1202020 1202012 1202011 1202010 1202002 1202001 1202000 1201222 1201221 1201220 1201212 1201211 1201210 1201202 1201201 1201200 1201122 1201121 1201120 1201112 1201111 1201110 1201102 1201101 1201100 1201022 1201021 1201020 1201012 1201011 1201010 1201002 1201001 1201000 1200222 1200221 1200220 1200212 1200211 1200210 1200210 1200201 1200200 1200122 1200121 1200120 1200112 1200111 1200110 1200102 1200101 1200100 1200022 1200021 1200020 1200012 1200011 1200010 1200011 1200010 1200001 1200000 1122222 1122221 1122220 1122212 1122211 1122210 1122202 1122201 1122200 1122122 1122121 1122120 1122112 1122111 1122110 1122102 1122101 1122100 1122022 1122021 1122020 1122012 1122011 1122010 1122002 1122001 1122000 1121000 1121000 1120222 1120221 1120220 1120212 1120211 1120210 1120202 1120201 1120200 1120122 1120121 1120120 1120112 1120111 1120110 1120102 1120101 1120100 1120022 1120021 1120020 1120012 1120011 1120010 1120002 1120001 1120000 1112222 1112221 1112220 1112212 1112211 1112210 1112202 1112201 1112200 1112122 1112121 1112120 1112112 1112111 1112110 1112102 1112101 1112101 1112102 1112101 1112100 1112022 1112021 1112020 1112012 1112011 1112010 1112002 1112001 1112000 1111222 1111221 1111220 1111212 1111211 1111210 1111202 1111201 1111200 1111122 1111121 1111120 1111112 1111111 1111110 1111102 1111101 1111100 1111022 1111021 1111020 1111012 1111011 1111010 1111002 1111001 1111000 1110222 1110221 1110220 1110212 1110211 1110210 1110202 1110201 1110200 1110122 1110121 1110120 1110112 1110111 1110110 1110102 1110101 1110100 1110012 1110011 1110010 1110002 1110001 1110000 1102222 1102221 1102220 1102212 1102211 1102210 1102202 1102201 1102200 1102122 1102121 1102120 1102112 1102111 1102110 1102102 1102101 1102100 1102012 1102011 1102010 1102002 1102001 1102000 1101222 1101221 1101220 1101212 1101211 1101210 1101202 1101201 1101200 1101122 1101121 1101120 1101112 1101111 1101110 1101102 1101101 1101100 1101022 1101021 1101020 1101012 1101011 1101010 1101002 1101000 1100222 1100221 1100220 1100212 1100211 1100210 1010202 1100202 1100201 1100200 1100122 1100121 1100120 1100112 1100111 1100110 1100102 1100101 1100100 1100022 1100021 1100020 1100012 1100011 1100010 1100002 1100001 1100000 1022222 1022221 1022220 1022212 1022211 1022210 1022202 1022201 1022200 1022122 1022121 1022120 1022112 1022111 1022110 1022102 1022101 1022100 1022022 1022021 1022020 1022012 1022011 1022012 1022010 1022002 1022001 1022000 1021222 1021221 1021220 1021212 1021211 1021210 1021202 1021201 1021200 1021122 1021121 1021120 1021112 1021111 1021110 1021102 1021101 1021100 1021022 1021021 1021020 1021001 1021000 1020122 1020121 1020120 1020112 1020111 1020110 1020102 1020101 1020100 1020022 1020021 1020020 1020012 1020011 1020010 1020010 1020002 1020001 1020000 1012222 1012221 1012220 1012212 1012211 1012210 1012202 1012201 1012200 1012122 1012121 1012120 1012112 1012112 1012111 1012110 1012102 1012101 1012100 1012022 1012021 1012020 1012012 1012011 1012010 1012002 1012001 1012000 1011222 1011221 1011220 1011212 1011211 1011210 1011202 1011201 1011200 1011122 1011121 1011120 1011112 1011111 1011110 1011102 1011101 1011100 1011022 1011021 1011020 1011012 1011011 1011010 1011002 1011001 1011000 1010222 1010221 1010220 1010212 1010211 1010210 1010202 1010201 1010200 1010122 1010121 1010122 1010120 1010121 1010111 1010111 1010102 1010101 1010100 1010022 1010021 1010020 1010012 1010011 1010010 1010002 1010001 1010000 1002222 1002221 1002220 1002212 1002211 1002210 1002202 1002201 1002200 1002122 1002121 1002120 1002112 1002111 1002110 1002102 1002101 1002100 1002022 1002121 1002120 1002112 1002111 1002110 1002102 1002101 1002100 1002022 1002021 1002020 1002012 1002011 1002010 1002002 1002001 1002000 1001222 1001221 1001220 1001212 1001211 1001210 1001202 1001201 1001200 1001122 1001121 1001120 1001120 1001111 1001110 1001102 1001101 1001100 1001022 1001021 1001020 1001012 1001011 1001010 1001002 1001001 1001000 1000222 1000221 1000220 1000212 1000211 1000201 1000200 1000122 1000121 1000120 1000112 1000111 1000110 1000102 1000100 1000022 1000021 1000020 1000012 1000011 1000010 1000002 1000001 1000000 222222 222221 222220 222212 222211 222210 222202 222201 222200 222022 222021 222020 222012 222011 222010 222002 222001 222000 221222 221221 222120 222112 222111 222110 222102 222101 222100 222022 222021 222020 222012 222011 222010 222002 222001 222000 221222 221221 221220 221212 221211 221210 221202 221201 221200 221122 221121 221120 221112 221111 221110 221102 221101 221102 221100 221022 221021 221020 221012 221011 221010 221002 221001 221000 220222 220221 220220 220212 220211 220210 220202 220201 220200 220122 220121 220120 220112 220111 220110 220102 220101 220100 220022 220021 220020 220012 220011 220010 220002 220001 220000 212222 212221 212220 212212 212211 212210 212202 212201 212200 212122 212121 212120 212112 212112 212111 212110 212102 212101 212100 212022 212021 212020 212012 212011 212010 221201 212001 212000 211222 211221 211220 211212 211211 211210 211202 211201 211202 211210 211201 211200 211122 211121 211120 211112 211111 211110 211102 211101 211100 211022 211021 211020 211012 211011 211012 211011 211010 211002 211001 211000 210222 210221 210220 210212 210211 210210 210202 210200 201000 200222 200221 200220 200212 200211 200210 200202 200201 200200 200122 200121 200120 200112 200111 200110 200102 200101 200100 200022 200021 200020 200012 200011 200010 200002 200001 200000 122222 122221 122220 122202 122201 122200 122122 122121 122120 122112 122111 122110 122102 122101 122100 122022 122021 122020 122002 122001 122000 121222 121220 121201 121200 121122 121121 121120 121112 121111 121110 121102 121101 121102 121101 121100 121022 121021 121020 121012 121011 121010 121002 121000 120222 120221 120220 120212 120211 120210 120202 120201 120200 120122 120121 120120 120112 120111 120110 120120 120112 120111 120110 120102 120101 120100 102222 120200 120122 120121 120120 120112 120111 120110 120102 120101 120100 120022 120021 120020 120012 120011 120010 120002 120001 120000 112222 112221 112220 112212 112211 112210 112202 112201 112200 112122 112121 112120 112112 112111 112110 112102 112101 112100 112022 112021 112020 112012 112011 112010 112002 112001 112000 111222 111221 111220 111212 111211 111210 111202 111201 111200 111122 111121 111120 111112 111111 111110 111102 111101 111100 111022 111021 111020 111012 111011 111010 111002 111001 111000 110222 110221 110220 110221 110220 110211 110210 110202 110201 110200 110122 110121 110120 110112 110111 110110 110102 110101 110101 110100 110022 110021 110020 110012 110011 110010 110002 110001 110000 102222 102221 102220 102212 102211 102210 102202 102201 102200 102122 102121 102102 102101 102100 102022 102021 102020 102012 102011 102010 102002 102001 102000 101222 101221 101220 101212 101211 101201 101210 101201 101200 101122 101121 101120 101112 101111 101110 101102 101101 101100 101022 101021 101020 101011 101010 101002 101001 101000 100222 100221 100220 100212 100211 100201 100202 100201 100200 100122 100121 100120 100112 100111 100110 100102 100101 100100 100022 100021 100020 100012 100011 100010 100002 100001 100000 22222 22221 22220 22212 22211 22210 22202 22201 22200 22122 22112 22020 22020 22012 22011 22010 22002 22001 22000 21222 21221 21220 21212 21211 21210 21202 21201 21200 21122 21121 21120 21112 21111 21112 21111 21110 21102 21101 21100 21022 21021 21020 21012 21011 21010 21002 21001 21000 20222 20221 20220 20212 20211 20210 20202 20201 20202 20200 20122 20121 20120 20112 20111 20110 20102 20101 20100 20022 20021 20020 20012 20011 20010 20002 20001 20000 12222 12221 12220 12212 12211 12210 12202 12201 12200 12122 12121 12120 12112 12111 12110 12102 12101 12100 12022 12021 12020 12012 12011 12010 12002 12001 12000 11222 11221 11220 11212 11210 11202 11201 11202 11201 11200 11122 11121 11120 11112 11111 11110 11102 11101 11100 11022 11021 11020 11012 11011 11010 11002 11001 11000 10222 10220 10202 10200 10122 10121 10120 10112 10111 10110 10102 10101 10101 10100 10022 10020 10012 10011 10010 10002 10002 10001 10000 2222 2221 2220 2212 2211 2210 2202 2201 2200 2122 2121 2120 2112 2111 2110 2102 2101 2100 2022 2021 2012 2011 2010 2002 2001 2000 1222 1221 1220 1212 1211 1210 1202 1201 1200 1122 1121 1120 1112 1111 1110 1102 1101 1100 1022 1021 1020 1012 1011 1010 1002 1001 1000 222 221 220 212 211 210 202 201 200 112 111 110 102 101 100 22 21 20 12 11 10 2 1 0 1 2 3 10 11 12 13 20 21 22 3 30 31 31 33 100 103 110 113 120 123 130 133 200 203 210 211 213 220 223 230 231 233 300 303 301 302 303 313 320 323 330 331 332 333 10000 10003 10010 10013 10020 10023 10030 10033 10100 10103 10110 10113 10120 10230 10231 10232 10233 10300 10303 10310 10313 10320 10323 10330 10331 10332 10333 11000 11001 11003 11010 11011 11012 11013 11020 11023 11030 11031 11032 11033 11100 11103 11110 11111 11113 11120 11130 11131 11132 11133 11200 11203 11213 11220 11223 11230 11233 11300 11303 11313 11323 11330 13333 20000 20001 20002 20003 20010 20011 20012 20013 20020 20021 20022 20023 20030 20031 20032 20033 20100 20101 20103 20110 20111 20113 20120 20113 20112 20111 20110 20103 20102 20101 20100 20033 20032 20031 20030 20030 20022 20021 20020 20013 20012 20011 20010 20003 20002 20001 20000 13333 13332 13331 13330 13323 13322 13321 13320 13313 13312 13311 13310 13303 13302 13301 13300 13233 13232 13231 13230 13223 13222 13221 13220 13213 13212 13211 13210 13203 13202 13201 13200 13133 13132 13131 13130 13123 13122 13121 13120 13113 13112 13111 13110 13103 13102 13101 13100 13033 13032 13031 13030 13023 13022 13021 13020 13013 13011 13010 13003 13002 13001 13000 12333 12332 12331 12330 12323 12322 12321 12320 12313 12312 12311 12310 12303 12302 12301 12300 12233 12232 12231 12230 12223 12222 12221 12220 12213 12211 12212 12210 12203 12202 12201 12200 12133 12132 12131 12130 12123 12122 12121 12120 12113 12112 12111 12110 12103 12102 12101 12100 12033 12032 12031 12030 12023 12001 12000 11333 11332 11331 11330 11323 11322 11321 11320 11313 11312 11311 11310 11303 11302 11301 11300 11233 11232 11231 11230 11223 11222 11221 11220 11213 11212 11211 11203 11202 11201 11200 11133 11132 11131 11130 11122 11121 11120 11113 11112 11111 11110 11103 11102 11101 11100 11033 11032 11013 11012 11011 11010 11003 11002 11001 11000 10333 10332 10331 10330 10323 10322 10321 10320 10313 10312 10311 10310 10303 10301 10300 10233 10232 10231 10230 10223 10222 10221 10220 10213 10212 10211 10210 10203 10202 10201 12000 10200 10133 10132 10131 10130 10123 10122 10121 10120 10113 10112 10111 10110 10103 10102 10101 10100 10033 10032 10031 10030 10023 10022 10021 10020 10013 10012 10011 10010 10003 10002 10001 10000 3333 3332 3331 3330 3323 3322 3321 3320 3313 3312 3311 3310 3303 3302 3301 3300 2333 2332 2331 2330 2323 2322 2321 2320 2313 2311 2310 2303 2302 2301 2300 2233 2230 2223 2222 2221 2220 2213 2212 2211 2210 2203 2202 2201 2200 2133 2132 2131 2130 2123 2122 2121 2120 2113 2112 2111 2110 2103 2102 2101 2100 2033 2032 2031 2030 2023 2022 2021 2020 2013 2012 2011 2010 2003 2002 2001 2000 1333 1332 1331 1330 1323 1322 1321 1320 1313 1312 1311 1310 1303 1302 1301 1300 1233 1232 1231 1230 1223 1222 1221 1220 1213 1212 1211 1210 1203 1202 1201 1200 1133 1132 1131 1130 1123 1122 1121 1120 1113 1112 1111 1110 1103 1102 1101 1100 1033 1032 1031 1030 1023 1022 1021 1020 1013 1012 1011 1010 1003 1002 1010 1001 1000 333 332 331 330 323 322 321 320 313 312 311 310 303 302 301 300 233 232 231 230 223 222 221 220 213 212 211 210 203 202 201 200 133 132 131 130 123 122 121 120 113 112 111 101 100 33 32 31 30 23 22 21 20 13 12 11 10 3 2 1 01 1