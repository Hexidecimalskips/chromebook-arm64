2 10 11 12 20 21 22 100 101 102 110 111 112 120 121 122 200 210 211 212 220 221 222 1000 1001 1002 1010 1011 1012 1020 1021 1022 1100 1101 1102 1110 1111 1112 1120 1121 1122 1200 1201 1202 1210 1211 1212 1220 1221 1222 2000 2001 2002 2010 2011 2102 2020 2021 2022 2100 2101 2102 2110 2111 2112 2120 2121 2122 2200 2201 2202 2210 2211 2212 2220 2221 2222 10000 10001 10002 10010 10011 10012 10020 10021 10022 10100 10101 10102 10110 10111 10112 10120 10121 10122 10200 10201 10202 10210 10211 10212 10220 10211 10221 10222 11000 11001 11002 11010 11011 11012 11020 11021 11022 11100 11101 11102 11110 11111 11112 11120 11121 11122 11200 11201 11202 11210 11211 11212 11220 11221 11222 12000 12001 12002 12010 12011 12012 12020 12021 12022 12100 12101 12102 12110 12111 12112 12120 1221 12122 12200 12201 12202 20000 12210 12211 12212 12220 12221 12222 20000 20001 20002 20010 20011 20012 20020 20021 20022 20100 20101 20102 20110 20111 20112 20120 20121 20122 20200 20201 20202 20201 20212 20220 20221 20222 21000 21001 21002 21010 21011 21012 21020 2021 21022 21100 2110 21102 21110 21111 21112 21120 21121 21212 21200 21201 21202 21210 21211 21212 21220 21221 21222 22000 22001 22200 22201 22202 22210 22211 22212 22220 22221 22222 1000000 100001 100002 100010 100011 100012 100020 100021 100022 100100 100101 100102 100110 100111 100112 100120 100121 100122 100200 100201 100202 100210 100211 100212 100220 100221 100222 101000 101001 101002 101010 101011 101012 101020 101021 101022 101100 101101 101102 101110 101111 101112 101120 101121 01112 101122 101200 101201 101202 101210 101211 101212 101220 101221 101222 102000 102001 102002 102010 102011 102012 102020 102021 102022 102100 102101 102102 102110 102111 102112 102120 102121 102122 102200 102201 102202 102210 102211 102212 102220 102221 102222 110000 110001 110002 110010 110011 110012 110021 110022 110100 110101 110102 110110 110111 110112 110120 110121 110122 110200 110202 110210 110211 110212 110220 110221 110222 111000 111001 111002 111010 111011 111012 111020 111021 111022 111100 111101 111102 111110 111111 111112 111120 111200 111201 111202 111210 111211 111212 111220 111221 111222 112000 112001 112002 112200 112201 112202 112210 112211 112212 112220 112221 112222 120000 120001 120002 120010 122000 122001 122002 122010 122011 122012 122020 122021 122022 122100 122102 122110 122111 122112 122120 122121 122122 122200 122201 122202 122210 122211 122212 122220 122221 122222 200000 200002 200010 200011 200012 200020 200021 200022 200100 200101 200102 200110 200111 200112 200120 200121 200122 200200 200201 200202 200210 200211 200212 200220 200221 200222 201000 201001 201002 201010 201011 201012 201020 201021 201022 201100 201101 201102 201110 201111 201112 201120 201121 201122 201200 201201 201202 201210 201211 201212 201220 201221 201222 202000 202001 202002 202010 2020211 202012 202020 202021 202022 202100 202101 0