100010000 1 10 11 100 101 110 111 1000 1001 1010 1011 1100 1101 1110 1111 10000 10001 10010 10011 10100 10101 10110 10111 11000 11001 11010 11011 11100 11101 11110 11111 100000 100001 100010 100011 100100 100101 100110 100111 101000 101001 101010 101011 101100 101101 101110 101111 110000 110001 110010 110011 110100 110101 110110 110111 111000 111001 111010 111011 111100 111101 111110 111111 1000000 10001000 10001001 10001010 10001011 10001100 1001101 10001101 10001110 10001111 10010000 10010001 10100010 10010011 10011000 10010101 10010110 10010111 10011000 10011001 10011010 10011011 10011100 10011101 10011110 10011111 10100000 10100001 10100010 10100011 10100100 10100101 10100110 10100111 10101000 10101001 10101011 10101100 10101111 10110000 10110001 10111100 10111101 10111110 10111111 11000000 11100000 11100001 11100010 11100011 11100100 11100101 11100110 11100111 11101000 11101001 11101010 11101011 11101100 11101101 11101110 11101111 11110000 11110001 11110010 11110011 11110100 11110101 11110110 11110111 11111000 11111001 11111010 11111101 11111110 11111111 11111110 11111101 11111100 11111011 11111010 11111001 11111000 11110111 11110110 11110101 11110100 11110011 11110010 11110001 11110000 11110111 11011111 11011110 11011101 11011100 11011011 11011010 11011001 11011000 11010111 11010110 11010101 11010100 11010011 11010010 11010001 11010000 11010000 11001111 11001110 11001010 11000111 11000110 11000101 11000100 11000010 11000001 11000000 10111111 10111110 10011111 10011110 10001111 10001110 10001101 10001100 10001011 10001010 10001001 10001000 10000111 10000101 10000100 10000011 10000010 10000001 10000000 01111111 00111111 00111110 00011111 00011110 00001111 00001110 00000111 00000110 00000010 00000000 1